library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity TEST is
  port (
    CLK      : in std_logic; -- 50 MHz system clock
    NRST     : in std_logic; -- Active-low asynchronous reset
    ADC_CSN  : out std_logic; -- ADC SPI chip-select
    ADC_SCLK : out std_logic; -- ADC SPI SCLK
    ADC_MOSI : out std_logic; -- ADC SPI MOSI
    ADC_MISO : in std_logic;  -- ADC SPI MISO
    LEDS     : out std_logic_vector(7 downto 0) -- 8-bit ADC OUTPUT
  );
end TEST;

architecture behavioral of TEST is

  constant SPI_CLK_DIV : integer := 25;
  constant DATA_WIDTH  : integer := 16; -- for ADC128S022

  type state_type is (ST_IDLE, ST_START, ST_SCK_H, ST_SCK_L, ST_WAIT);
  signal state : state_type := ST_IDLE;

  signal cs_n : std_logic := '1';
  signal sclk : std_logic := '0';
  signal mosi : std_logic := '0';

  signal bit_index : integer range 0 to DATA_WIDTH - 1 := 0;
  signal adc_data  : std_logic_vector(11 downto 0)  := (others => '0');
  signal channel   : std_logic_vector(2 downto 0)   := "111";

  signal shift_en  : std_logic := '0';
  signal shift_reg : std_logic_vector(DATA_WIDTH - 1 downto 0);

  constant WAIT_CNT_MAX : integer := 31;
  signal wait_cnt       : integer := 0;

begin

  adc_csn  <= cs_n;
  adc_sclk <= sclk;
  adc_mosi <= mosi;

  --LEDS <= adc_data(11 downto 4); -- show 8-bit ADC value directly to LEDs

  process (adc_data)
    variable leds_on : integer range 0 to 7;
    variable value   : integer range 0 to 255;
  begin
    value   := to_integer(unsigned(adc_data(11 downto 4)));
    value   := value / 32;
    leds_on := value;
    LEDS <= (others => '0'); -- Default to all LEDs OFF
    LEDS(leds_on downto 0) <= (others => '1'); -- Turn ON the corresponding LEDs
  end process;

  process (CLK, NRST)
    variable count : integer range 0 to SPI_CLK_DIV - 1 := 0;
  begin
    if NRST = '0' then
      count := 0;
      shift_en <= '0';
    elsif rising_edge(CLK) then
      if count = SPI_CLK_DIV - 1 then
        count := 0;
        shift_en <= '1';
      else
        count := count + 1;
        shift_en <= '0';
      end if;
    end if;
  end process;

  process (CLK, NRST)
  begin
    if NRST = '0' then
      cs_n      <= '1';
      mosi      <= '0';
      sclk      <= '0';
      adc_data  <= (others => '0');
      channel   <= (others => '0');
      bit_index <= 0;
      wait_cnt  <= 0;
      state     <= ST_IDLE;

    elsif rising_edge(CLK) then

      case state is
        when ST_IDLE =>
          bit_index <= 0;
          channel   <= "111"; -- Select channel ADC_IN1
          cs_n      <= '1';
          sclk      <= '1';
          state     <= ST_START;

        when ST_START  =>
          shift_reg  <= (others => '0');
          shift_reg(13 downto 11) <= channel; -- for ADC128S022
          cs_n   <= '0';
          state  <= ST_SCK_L;

        when ST_SCK_L =>
          if shift_en = '1' then
            sclk  <= '0';
            mosi  <= shift_reg(shift_reg'left);
            state <= ST_SCK_H;
          end if;

        when ST_SCK_H =>
          if shift_en = '1' then
            sclk      <= '1';
            shift_reg <= shift_reg(shift_reg'left - 1 downto 0) & adc_miso;
            if bit_index = DATA_WIDTH - 1 then
              cs_n     <= '1';
              wait_cnt <= WAIT_CNT_MAX;
              state    <= ST_WAIT;
            else
              bit_index <= bit_index + 1;
              state     <= ST_SCK_L;
            end if;
          end if;

        when ST_WAIT =>
          adc_data <= shift_reg(11 downto 0);
          if wait_cnt = 0 then
            state <= ST_IDLE;
          else
            wait_cnt <= wait_cnt - 1;
          end if;

        when others =>
          state <= ST_IDLE;
      end case;
    end if;
  end process;

end behavioral;